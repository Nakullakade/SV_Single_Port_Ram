class configuration;
  virtual s_interface vif;
  mailbox gen2Driv;
  mailbox ip_mon2scbd;
  mailbox op_mon2scbd;
  mailbox ip_mon2conv;
  mailbox op_mon2conv;
endclass