package s_package;
`include "define.sv"
`include "packet.sv"
`include "configuration.sv"
`include "Scoreboard.sv"
`include "coverage_collector.sv"
`include "op_monitor.sv"
`include "ip_monitor.sv"
`include "Driver.sv"
`include "generator.sv"
`include "environment.sv"
`include "test.sv"
endpackage