typedef virtual s_interface.tb intf_t1;
